/********|********|********|********|********|********|********|********/
/*                        TRABALHO IV SD                               */
/* File:   fpu_types.sv                                                */
/* Author: Fernando Acauan                                             */
/*                                                                     */
/********|********|********|********|********|********|********|********/
/********|********|********|********|********|********|********|********/

/********|********|********|********|********|********|********|********/
/*                                                                     */
/*                           FPU_types                                 */
/*                                                                     */
/********|********|********|********|********|********|********|********/

package FPU_types;

    typedef enum logic [3:0] { EXACT, OVERFLOW, UNDERFLOW, INEXACT } g_eStatus;

endpackage

/********|********|********|********|********|********|********|********/

